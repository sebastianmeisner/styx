----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:00:49 05/21/2013 
-- Design Name: 
-- Module Name:    test_circuit - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity InverterChain is
	generic (
		n: positive range 2 to 16384 := 1024
	);
	port ( 	
		clk : in std_logic; 
		rst : in std_logic;
		intr_out : out std_logic_vector(127 downto 0)
	);
end InverterChain;

architecture structural of InverterChain is 
	-- Interne Signale
	-- Verbindungen zwischen den einzelnen Inverter-FlipFlop Elementen
	-- intern-Signale verbindet alle Elemente untereinander
	-- intern_se verbindet Start- mit End-Element
	signal intern : std_logic_vector(1 to n-1);
	signal intern_se : std_logic;
	signal reset : std_logic;
	
	signal a : std_logic := '0';
	signal b : std_logic := '0';
	
	-- keep-Attribut zur Vermeidung der Wegoptimierung durch
	-- Synthese Werkzeug
	attribute keep : string;
	attribute keep of intern : signal is "true";
	attribute keep of intern_se : signal is "true";
	
component InverterElemP 
	port (
		d : in  std_logic;
      clk : in  std_logic;
      q : out  std_logic;
		reset : in std_logic
	) ;
end component;

begin 

	-- Instanziieren der Inverter-Elemente
	-- und Verbinden der Elemente untereinander
	reg : for i in n downto 1 generate
		
		-- Betrachtung des ERSTEN Elements
		reg_begin: if i = 1 generate 
			InverterElem_begin: InverterElemP 
				port map (intern_se, clk, intern(i), reset) ;
		end generate ;

		-- Betrachtung der MITTLEREN Elemente
		reg_middle_p: if i > 1 and i < n generate 
			InverterElem_middle_p: InverterElemP 
				port map (intern(i-1), clk, intern(i), reset) ;
		end generate ;

		-- Betrachtung des LETZTEN Elements
		reg_end: if i = n generate 
			InverterElem_end: InverterElemP 
				port map (intern(i-1), clk, intern_se, reset) ;
		end generate ;
	end generate ;
	
	
	process(clk, rst)
	begin
		if(rst = '1') then
			intr_out(0) 	 <= 	 '0';--(intern(1) AND intern(2) AND intern(3) AND intern(4) AND intern(5) AND intern(6) AND intern(7) AND intern(8)) OR ((NOT intern(1)) AND (NOT intern(2)) AND (NOT intern(3)) AND (NOT intern(4)) AND (NOT intern(5)) AND (NOT intern(6)) AND (NOT intern(7)) AND (NOT intern(8)));
			intr_out(1) 	 <= 	 '0';--(intern(9) AND intern(10) AND intern(11) AND intern(12) AND intern(13) AND intern(14) AND intern(15) AND intern(16)) OR ((NOT intern(9)) AND (NOT intern(10)) AND (NOT intern(11)) AND (NOT intern(12)) AND (NOT intern(13)) AND (NOT intern(14)) AND (NOT intern(15)) AND (NOT intern(16)));
		elsif(clk = '1' and clk'event) then
			intr_out(0) 	 <= 	 intern(513);--(intern(1) AND intern(2) AND intern(3) AND intern(4) AND intern(5) AND intern(6) AND intern(7) AND intern(8)) OR ((NOT intern(1)) AND (NOT intern(2)) AND (NOT intern(3)) AND (NOT intern(4)) AND (NOT intern(5)) AND (NOT intern(6)) AND (NOT intern(7)) AND (NOT intern(8)));
			intr_out(1) 	 <= 	 intern(514);--(intern(9) AND intern(10) AND intern(11) AND intern(12) AND intern(13) AND intern(14) AND intern(15) AND intern(16)) OR ((NOT intern(9)) AND (NOT intern(10)) AND (NOT intern(11)) AND (NOT intern(12)) AND (NOT intern(13)) AND (NOT intern(14)) AND (NOT intern(15)) AND (NOT intern(16)));

		end if;
	end process;

--	intr_out(0) 	 <= 	 intern(513);--(intern(1) AND intern(2) AND intern(3) AND intern(4) AND intern(5) AND intern(6) AND intern(7) AND intern(8)) OR ((NOT intern(1)) AND (NOT intern(2)) AND (NOT intern(3)) AND (NOT intern(4)) AND (NOT intern(5)) AND (NOT intern(6)) AND (NOT intern(7)) AND (NOT intern(8)));
--	intr_out(1) 	 <= 	 intern(514);--(intern(9) AND intern(10) AND intern(11) AND intern(12) AND intern(13) AND intern(14) AND intern(15) AND intern(16)) OR ((NOT intern(9)) AND (NOT intern(10)) AND (NOT intern(11)) AND (NOT intern(12)) AND (NOT intern(13)) AND (NOT intern(14)) AND (NOT intern(15)) AND (NOT intern(16)));
--	intr_out(2) 	 <= 	 (intern(17) AND intern(18) AND intern(19) AND intern(20) AND intern(21) AND intern(22) AND intern(23) AND intern(24)) OR ((NOT intern(17)) AND (NOT intern(18)) AND (NOT intern(19)) AND (NOT intern(20)) AND (NOT intern(21)) AND (NOT intern(22)) AND (NOT intern(23)) AND (NOT intern(24)));
--	intr_out(3) 	 <= 	 (intern(25) AND intern(26) AND intern(27) AND intern(28) AND intern(29) AND intern(30) AND intern(31) AND intern(32)) OR ((NOT intern(25)) AND (NOT intern(26)) AND (NOT intern(27)) AND (NOT intern(28)) AND (NOT intern(29)) AND (NOT intern(30)) AND (NOT intern(31)) AND (NOT intern(32)));
--	intr_out(4) 	 <= 	 (intern(33) AND intern(34) AND intern(35) AND intern(36) AND intern(37) AND intern(38) AND intern(39) AND intern(40)) OR ((NOT intern(33)) AND (NOT intern(34)) AND (NOT intern(35)) AND (NOT intern(36)) AND (NOT intern(37)) AND (NOT intern(38)) AND (NOT intern(39)) AND (NOT intern(40)));
--	intr_out(5) 	 <= 	 (intern(41) AND intern(42) AND intern(43) AND intern(44) AND intern(45) AND intern(46) AND intern(47) AND intern(48)) OR ((NOT intern(41)) AND (NOT intern(42)) AND (NOT intern(43)) AND (NOT intern(44)) AND (NOT intern(45)) AND (NOT intern(46)) AND (NOT intern(47)) AND (NOT intern(48)));
--	intr_out(6) 	 <= 	 (intern(49) AND intern(50) AND intern(51) AND intern(52) AND intern(53) AND intern(54) AND intern(55) AND intern(56)) OR ((NOT intern(49)) AND (NOT intern(50)) AND (NOT intern(51)) AND (NOT intern(52)) AND (NOT intern(53)) AND (NOT intern(54)) AND (NOT intern(55)) AND (NOT intern(56)));
--	intr_out(7) 	 <= 	 (intern(57) AND intern(58) AND intern(59) AND intern(60) AND intern(61) AND intern(62) AND intern(63) AND intern(64)) OR ((NOT intern(57)) AND (NOT intern(58)) AND (NOT intern(59)) AND (NOT intern(60)) AND (NOT intern(61)) AND (NOT intern(62)) AND (NOT intern(63)) AND (NOT intern(64)));
--	intr_out(8) 	 <= 	 (intern(65) AND intern(66) AND intern(67) AND intern(68) AND intern(69) AND intern(70) AND intern(71) AND intern(72)) OR ((NOT intern(65)) AND (NOT intern(66)) AND (NOT intern(67)) AND (NOT intern(68)) AND (NOT intern(69)) AND (NOT intern(70)) AND (NOT intern(71)) AND (NOT intern(72)));
--	intr_out(9) 	 <= 	 (intern(73) AND intern(74) AND intern(75) AND intern(76) AND intern(77) AND intern(78) AND intern(79) AND intern(80)) OR ((NOT intern(73)) AND (NOT intern(74)) AND (NOT intern(75)) AND (NOT intern(76)) AND (NOT intern(77)) AND (NOT intern(78)) AND (NOT intern(79)) AND (NOT intern(80)));
--	intr_out(10) 	 <= 	 (intern(81) AND intern(82) AND intern(83) AND intern(84) AND intern(85) AND intern(86) AND intern(87) AND intern(88)) OR ((NOT intern(81)) AND (NOT intern(82)) AND (NOT intern(83)) AND (NOT intern(84)) AND (NOT intern(85)) AND (NOT intern(86)) AND (NOT intern(87)) AND (NOT intern(88)));
--	intr_out(11) 	 <= 	 (intern(89) AND intern(90) AND intern(91) AND intern(92) AND intern(93) AND intern(94) AND intern(95) AND intern(96)) OR ((NOT intern(89)) AND (NOT intern(90)) AND (NOT intern(91)) AND (NOT intern(92)) AND (NOT intern(93)) AND (NOT intern(94)) AND (NOT intern(95)) AND (NOT intern(96)));
--	intr_out(12) 	 <= 	 (intern(97) AND intern(98) AND intern(99) AND intern(100) AND intern(101) AND intern(102) AND intern(103) AND intern(104)) OR ((NOT intern(97)) AND (NOT intern(98)) AND (NOT intern(99)) AND (NOT intern(100)) AND (NOT intern(101)) AND (NOT intern(102)) AND (NOT intern(103)) AND (NOT intern(104)));
--	intr_out(13) 	 <= 	 (intern(105) AND intern(106) AND intern(107) AND intern(108) AND intern(109) AND intern(110) AND intern(111) AND intern(112)) OR ((NOT intern(105)) AND (NOT intern(106)) AND (NOT intern(107)) AND (NOT intern(108)) AND (NOT intern(109)) AND (NOT intern(110)) AND (NOT intern(111)) AND (NOT intern(112)));
--	intr_out(14) 	 <= 	 (intern(113) AND intern(114) AND intern(115) AND intern(116) AND intern(117) AND intern(118) AND intern(119) AND intern(120)) OR ((NOT intern(113)) AND (NOT intern(114)) AND (NOT intern(115)) AND (NOT intern(116)) AND (NOT intern(117)) AND (NOT intern(118)) AND (NOT intern(119)) AND (NOT intern(120)));
--	intr_out(15) 	 <= 	 (intern(121) AND intern(122) AND intern(123) AND intern(124) AND intern(125) AND intern(126) AND intern(127) AND intern(128)) OR ((NOT intern(121)) AND (NOT intern(122)) AND (NOT intern(123)) AND (NOT intern(124)) AND (NOT intern(125)) AND (NOT intern(126)) AND (NOT intern(127)) AND (NOT intern(128)));
--	intr_out(16) 	 <= 	 (intern(129) AND intern(130) AND intern(131) AND intern(132) AND intern(133) AND intern(134) AND intern(135) AND intern(136)) OR ((NOT intern(129)) AND (NOT intern(130)) AND (NOT intern(131)) AND (NOT intern(132)) AND (NOT intern(133)) AND (NOT intern(134)) AND (NOT intern(135)) AND (NOT intern(136)));
--	intr_out(17) 	 <= 	 (intern(137) AND intern(138) AND intern(139) AND intern(140) AND intern(141) AND intern(142) AND intern(143) AND intern(144)) OR ((NOT intern(137)) AND (NOT intern(138)) AND (NOT intern(139)) AND (NOT intern(140)) AND (NOT intern(141)) AND (NOT intern(142)) AND (NOT intern(143)) AND (NOT intern(144)));
--	intr_out(18) 	 <= 	 (intern(145) AND intern(146) AND intern(147) AND intern(148) AND intern(149) AND intern(150) AND intern(151) AND intern(152)) OR ((NOT intern(145)) AND (NOT intern(146)) AND (NOT intern(147)) AND (NOT intern(148)) AND (NOT intern(149)) AND (NOT intern(150)) AND (NOT intern(151)) AND (NOT intern(152)));
--	intr_out(19) 	 <= 	 (intern(153) AND intern(154) AND intern(155) AND intern(156) AND intern(157) AND intern(158) AND intern(159) AND intern(160)) OR ((NOT intern(153)) AND (NOT intern(154)) AND (NOT intern(155)) AND (NOT intern(156)) AND (NOT intern(157)) AND (NOT intern(158)) AND (NOT intern(159)) AND (NOT intern(160)));
--	intr_out(20) 	 <= 	 (intern(161) AND intern(162) AND intern(163) AND intern(164) AND intern(165) AND intern(166) AND intern(167) AND intern(168)) OR ((NOT intern(161)) AND (NOT intern(162)) AND (NOT intern(163)) AND (NOT intern(164)) AND (NOT intern(165)) AND (NOT intern(166)) AND (NOT intern(167)) AND (NOT intern(168)));
--	intr_out(21) 	 <= 	 (intern(169) AND intern(170) AND intern(171) AND intern(172) AND intern(173) AND intern(174) AND intern(175) AND intern(176)) OR ((NOT intern(169)) AND (NOT intern(170)) AND (NOT intern(171)) AND (NOT intern(172)) AND (NOT intern(173)) AND (NOT intern(174)) AND (NOT intern(175)) AND (NOT intern(176)));
--	intr_out(22) 	 <= 	 (intern(177) AND intern(178) AND intern(179) AND intern(180) AND intern(181) AND intern(182) AND intern(183) AND intern(184)) OR ((NOT intern(177)) AND (NOT intern(178)) AND (NOT intern(179)) AND (NOT intern(180)) AND (NOT intern(181)) AND (NOT intern(182)) AND (NOT intern(183)) AND (NOT intern(184)));
--	intr_out(23) 	 <= 	 (intern(185) AND intern(186) AND intern(187) AND intern(188) AND intern(189) AND intern(190) AND intern(191) AND intern(192)) OR ((NOT intern(185)) AND (NOT intern(186)) AND (NOT intern(187)) AND (NOT intern(188)) AND (NOT intern(189)) AND (NOT intern(190)) AND (NOT intern(191)) AND (NOT intern(192)));
--	intr_out(24) 	 <= 	 (intern(193) AND intern(194) AND intern(195) AND intern(196) AND intern(197) AND intern(198) AND intern(199) AND intern(200)) OR ((NOT intern(193)) AND (NOT intern(194)) AND (NOT intern(195)) AND (NOT intern(196)) AND (NOT intern(197)) AND (NOT intern(198)) AND (NOT intern(199)) AND (NOT intern(200)));
--	intr_out(25) 	 <= 	 (intern(201) AND intern(202) AND intern(203) AND intern(204) AND intern(205) AND intern(206) AND intern(207) AND intern(208)) OR ((NOT intern(201)) AND (NOT intern(202)) AND (NOT intern(203)) AND (NOT intern(204)) AND (NOT intern(205)) AND (NOT intern(206)) AND (NOT intern(207)) AND (NOT intern(208)));
--	intr_out(26) 	 <= 	 (intern(209) AND intern(210) AND intern(211) AND intern(212) AND intern(213) AND intern(214) AND intern(215) AND intern(216)) OR ((NOT intern(209)) AND (NOT intern(210)) AND (NOT intern(211)) AND (NOT intern(212)) AND (NOT intern(213)) AND (NOT intern(214)) AND (NOT intern(215)) AND (NOT intern(216)));
--	intr_out(27) 	 <= 	 (intern(217) AND intern(218) AND intern(219) AND intern(220) AND intern(221) AND intern(222) AND intern(223) AND intern(224)) OR ((NOT intern(217)) AND (NOT intern(218)) AND (NOT intern(219)) AND (NOT intern(220)) AND (NOT intern(221)) AND (NOT intern(222)) AND (NOT intern(223)) AND (NOT intern(224)));
--	intr_out(28) 	 <= 	 (intern(225) AND intern(226) AND intern(227) AND intern(228) AND intern(229) AND intern(230) AND intern(231) AND intern(232)) OR ((NOT intern(225)) AND (NOT intern(226)) AND (NOT intern(227)) AND (NOT intern(228)) AND (NOT intern(229)) AND (NOT intern(230)) AND (NOT intern(231)) AND (NOT intern(232)));
--	intr_out(29) 	 <= 	 (intern(233) AND intern(234) AND intern(235) AND intern(236) AND intern(237) AND intern(238) AND intern(239) AND intern(240)) OR ((NOT intern(233)) AND (NOT intern(234)) AND (NOT intern(235)) AND (NOT intern(236)) AND (NOT intern(237)) AND (NOT intern(238)) AND (NOT intern(239)) AND (NOT intern(240)));
--	intr_out(30) 	 <= 	 (intern(241) AND intern(242) AND intern(243) AND intern(244) AND intern(245) AND intern(246) AND intern(247) AND intern(248)) OR ((NOT intern(241)) AND (NOT intern(242)) AND (NOT intern(243)) AND (NOT intern(244)) AND (NOT intern(245)) AND (NOT intern(246)) AND (NOT intern(247)) AND (NOT intern(248)));
--	intr_out(31) 	 <= 	 (intern(249) AND intern(250) AND intern(251) AND intern(252) AND intern(253) AND intern(254) AND intern(255) AND intern(256)) OR ((NOT intern(249)) AND (NOT intern(250)) AND (NOT intern(251)) AND (NOT intern(252)) AND (NOT intern(253)) AND (NOT intern(254)) AND (NOT intern(255)) AND (NOT intern(256)));
--	intr_out(32) 	 <= 	 (intern(257) AND intern(258) AND intern(259) AND intern(260) AND intern(261) AND intern(262) AND intern(263) AND intern(264)) OR ((NOT intern(257)) AND (NOT intern(258)) AND (NOT intern(259)) AND (NOT intern(260)) AND (NOT intern(261)) AND (NOT intern(262)) AND (NOT intern(263)) AND (NOT intern(264)));
--	intr_out(33) 	 <= 	 (intern(265) AND intern(266) AND intern(267) AND intern(268) AND intern(269) AND intern(270) AND intern(271) AND intern(272)) OR ((NOT intern(265)) AND (NOT intern(266)) AND (NOT intern(267)) AND (NOT intern(268)) AND (NOT intern(269)) AND (NOT intern(270)) AND (NOT intern(271)) AND (NOT intern(272)));
--	intr_out(34) 	 <= 	 (intern(273) AND intern(274) AND intern(275) AND intern(276) AND intern(277) AND intern(278) AND intern(279) AND intern(280)) OR ((NOT intern(273)) AND (NOT intern(274)) AND (NOT intern(275)) AND (NOT intern(276)) AND (NOT intern(277)) AND (NOT intern(278)) AND (NOT intern(279)) AND (NOT intern(280)));
--	intr_out(35) 	 <= 	 (intern(281) AND intern(282) AND intern(283) AND intern(284) AND intern(285) AND intern(286) AND intern(287) AND intern(288)) OR ((NOT intern(281)) AND (NOT intern(282)) AND (NOT intern(283)) AND (NOT intern(284)) AND (NOT intern(285)) AND (NOT intern(286)) AND (NOT intern(287)) AND (NOT intern(288)));
--	intr_out(36) 	 <= 	 (intern(289) AND intern(290) AND intern(291) AND intern(292) AND intern(293) AND intern(294) AND intern(295) AND intern(296)) OR ((NOT intern(289)) AND (NOT intern(290)) AND (NOT intern(291)) AND (NOT intern(292)) AND (NOT intern(293)) AND (NOT intern(294)) AND (NOT intern(295)) AND (NOT intern(296)));
--	intr_out(37) 	 <= 	 (intern(297) AND intern(298) AND intern(299) AND intern(300) AND intern(301) AND intern(302) AND intern(303) AND intern(304)) OR ((NOT intern(297)) AND (NOT intern(298)) AND (NOT intern(299)) AND (NOT intern(300)) AND (NOT intern(301)) AND (NOT intern(302)) AND (NOT intern(303)) AND (NOT intern(304)));
--	intr_out(38) 	 <= 	 (intern(305) AND intern(306) AND intern(307) AND intern(308) AND intern(309) AND intern(310) AND intern(311) AND intern(312)) OR ((NOT intern(305)) AND (NOT intern(306)) AND (NOT intern(307)) AND (NOT intern(308)) AND (NOT intern(309)) AND (NOT intern(310)) AND (NOT intern(311)) AND (NOT intern(312)));
--	intr_out(39) 	 <= 	 (intern(313) AND intern(314) AND intern(315) AND intern(316) AND intern(317) AND intern(318) AND intern(319) AND intern(320)) OR ((NOT intern(313)) AND (NOT intern(314)) AND (NOT intern(315)) AND (NOT intern(316)) AND (NOT intern(317)) AND (NOT intern(318)) AND (NOT intern(319)) AND (NOT intern(320)));
--	intr_out(40) 	 <= 	 (intern(321) AND intern(322) AND intern(323) AND intern(324) AND intern(325) AND intern(326) AND intern(327) AND intern(328)) OR ((NOT intern(321)) AND (NOT intern(322)) AND (NOT intern(323)) AND (NOT intern(324)) AND (NOT intern(325)) AND (NOT intern(326)) AND (NOT intern(327)) AND (NOT intern(328)));
--	intr_out(41) 	 <= 	 (intern(329) AND intern(330) AND intern(331) AND intern(332) AND intern(333) AND intern(334) AND intern(335) AND intern(336)) OR ((NOT intern(329)) AND (NOT intern(330)) AND (NOT intern(331)) AND (NOT intern(332)) AND (NOT intern(333)) AND (NOT intern(334)) AND (NOT intern(335)) AND (NOT intern(336)));
--	intr_out(42) 	 <= 	 (intern(337) AND intern(338) AND intern(339) AND intern(340) AND intern(341) AND intern(342) AND intern(343) AND intern(344)) OR ((NOT intern(337)) AND (NOT intern(338)) AND (NOT intern(339)) AND (NOT intern(340)) AND (NOT intern(341)) AND (NOT intern(342)) AND (NOT intern(343)) AND (NOT intern(344)));
--	intr_out(43) 	 <= 	 (intern(345) AND intern(346) AND intern(347) AND intern(348) AND intern(349) AND intern(350) AND intern(351) AND intern(352)) OR ((NOT intern(345)) AND (NOT intern(346)) AND (NOT intern(347)) AND (NOT intern(348)) AND (NOT intern(349)) AND (NOT intern(350)) AND (NOT intern(351)) AND (NOT intern(352)));
--	intr_out(44) 	 <= 	 (intern(353) AND intern(354) AND intern(355) AND intern(356) AND intern(357) AND intern(358) AND intern(359) AND intern(360)) OR ((NOT intern(353)) AND (NOT intern(354)) AND (NOT intern(355)) AND (NOT intern(356)) AND (NOT intern(357)) AND (NOT intern(358)) AND (NOT intern(359)) AND (NOT intern(360)));
--	intr_out(45) 	 <= 	 (intern(361) AND intern(362) AND intern(363) AND intern(364) AND intern(365) AND intern(366) AND intern(367) AND intern(368)) OR ((NOT intern(361)) AND (NOT intern(362)) AND (NOT intern(363)) AND (NOT intern(364)) AND (NOT intern(365)) AND (NOT intern(366)) AND (NOT intern(367)) AND (NOT intern(368)));
--	intr_out(46) 	 <= 	 (intern(369) AND intern(370) AND intern(371) AND intern(372) AND intern(373) AND intern(374) AND intern(375) AND intern(376)) OR ((NOT intern(369)) AND (NOT intern(370)) AND (NOT intern(371)) AND (NOT intern(372)) AND (NOT intern(373)) AND (NOT intern(374)) AND (NOT intern(375)) AND (NOT intern(376)));
--	intr_out(47) 	 <= 	 (intern(377) AND intern(378) AND intern(379) AND intern(380) AND intern(381) AND intern(382) AND intern(383) AND intern(384)) OR ((NOT intern(377)) AND (NOT intern(378)) AND (NOT intern(379)) AND (NOT intern(380)) AND (NOT intern(381)) AND (NOT intern(382)) AND (NOT intern(383)) AND (NOT intern(384)));
--	intr_out(48) 	 <= 	 (intern(385) AND intern(386) AND intern(387) AND intern(388) AND intern(389) AND intern(390) AND intern(391) AND intern(392)) OR ((NOT intern(385)) AND (NOT intern(386)) AND (NOT intern(387)) AND (NOT intern(388)) AND (NOT intern(389)) AND (NOT intern(390)) AND (NOT intern(391)) AND (NOT intern(392)));
--	intr_out(49) 	 <= 	 (intern(393) AND intern(394) AND intern(395) AND intern(396) AND intern(397) AND intern(398) AND intern(399) AND intern(400)) OR ((NOT intern(393)) AND (NOT intern(394)) AND (NOT intern(395)) AND (NOT intern(396)) AND (NOT intern(397)) AND (NOT intern(398)) AND (NOT intern(399)) AND (NOT intern(400)));
--	intr_out(50) 	 <= 	 (intern(401) AND intern(402) AND intern(403) AND intern(404) AND intern(405) AND intern(406) AND intern(407) AND intern(408)) OR ((NOT intern(401)) AND (NOT intern(402)) AND (NOT intern(403)) AND (NOT intern(404)) AND (NOT intern(405)) AND (NOT intern(406)) AND (NOT intern(407)) AND (NOT intern(408)));
--	intr_out(51) 	 <= 	 (intern(409) AND intern(410) AND intern(411) AND intern(412) AND intern(413) AND intern(414) AND intern(415) AND intern(416)) OR ((NOT intern(409)) AND (NOT intern(410)) AND (NOT intern(411)) AND (NOT intern(412)) AND (NOT intern(413)) AND (NOT intern(414)) AND (NOT intern(415)) AND (NOT intern(416)));
--	intr_out(52) 	 <= 	 (intern(417) AND intern(418) AND intern(419) AND intern(420) AND intern(421) AND intern(422) AND intern(423) AND intern(424)) OR ((NOT intern(417)) AND (NOT intern(418)) AND (NOT intern(419)) AND (NOT intern(420)) AND (NOT intern(421)) AND (NOT intern(422)) AND (NOT intern(423)) AND (NOT intern(424)));
--	intr_out(53) 	 <= 	 (intern(425) AND intern(426) AND intern(427) AND intern(428) AND intern(429) AND intern(430) AND intern(431) AND intern(432)) OR ((NOT intern(425)) AND (NOT intern(426)) AND (NOT intern(427)) AND (NOT intern(428)) AND (NOT intern(429)) AND (NOT intern(430)) AND (NOT intern(431)) AND (NOT intern(432)));
--	intr_out(54) 	 <= 	 (intern(433) AND intern(434) AND intern(435) AND intern(436) AND intern(437) AND intern(438) AND intern(439) AND intern(440)) OR ((NOT intern(433)) AND (NOT intern(434)) AND (NOT intern(435)) AND (NOT intern(436)) AND (NOT intern(437)) AND (NOT intern(438)) AND (NOT intern(439)) AND (NOT intern(440)));
--	intr_out(55) 	 <= 	 (intern(441) AND intern(442) AND intern(443) AND intern(444) AND intern(445) AND intern(446) AND intern(447) AND intern(448)) OR ((NOT intern(441)) AND (NOT intern(442)) AND (NOT intern(443)) AND (NOT intern(444)) AND (NOT intern(445)) AND (NOT intern(446)) AND (NOT intern(447)) AND (NOT intern(448)));
--	intr_out(56) 	 <= 	 (intern(449) AND intern(450) AND intern(451) AND intern(452) AND intern(453) AND intern(454) AND intern(455) AND intern(456)) OR ((NOT intern(449)) AND (NOT intern(450)) AND (NOT intern(451)) AND (NOT intern(452)) AND (NOT intern(453)) AND (NOT intern(454)) AND (NOT intern(455)) AND (NOT intern(456)));
--	intr_out(57) 	 <= 	 (intern(457) AND intern(458) AND intern(459) AND intern(460) AND intern(461) AND intern(462) AND intern(463) AND intern(464)) OR ((NOT intern(457)) AND (NOT intern(458)) AND (NOT intern(459)) AND (NOT intern(460)) AND (NOT intern(461)) AND (NOT intern(462)) AND (NOT intern(463)) AND (NOT intern(464)));
--	intr_out(58) 	 <= 	 (intern(465) AND intern(466) AND intern(467) AND intern(468) AND intern(469) AND intern(470) AND intern(471) AND intern(472)) OR ((NOT intern(465)) AND (NOT intern(466)) AND (NOT intern(467)) AND (NOT intern(468)) AND (NOT intern(469)) AND (NOT intern(470)) AND (NOT intern(471)) AND (NOT intern(472)));
--	intr_out(59) 	 <= 	 (intern(473) AND intern(474) AND intern(475) AND intern(476) AND intern(477) AND intern(478) AND intern(479) AND intern(480)) OR ((NOT intern(473)) AND (NOT intern(474)) AND (NOT intern(475)) AND (NOT intern(476)) AND (NOT intern(477)) AND (NOT intern(478)) AND (NOT intern(479)) AND (NOT intern(480)));
--	intr_out(60) 	 <= 	 (intern(481) AND intern(482) AND intern(483) AND intern(484) AND intern(485) AND intern(486) AND intern(487) AND intern(488)) OR ((NOT intern(481)) AND (NOT intern(482)) AND (NOT intern(483)) AND (NOT intern(484)) AND (NOT intern(485)) AND (NOT intern(486)) AND (NOT intern(487)) AND (NOT intern(488)));
--	intr_out(61) 	 <= 	 (intern(489) AND intern(490) AND intern(491) AND intern(492) AND intern(493) AND intern(494) AND intern(495) AND intern(496)) OR ((NOT intern(489)) AND (NOT intern(490)) AND (NOT intern(491)) AND (NOT intern(492)) AND (NOT intern(493)) AND (NOT intern(494)) AND (NOT intern(495)) AND (NOT intern(496)));
--	intr_out(62) 	 <= 	 (intern(497) AND intern(498) AND intern(499) AND intern(500) AND intern(501) AND intern(502) AND intern(503) AND intern(504)) OR ((NOT intern(497)) AND (NOT intern(498)) AND (NOT intern(499)) AND (NOT intern(500)) AND (NOT intern(501)) AND (NOT intern(502)) AND (NOT intern(503)) AND (NOT intern(504)));
--	intr_out(63) 	 <= 	 (intern(505) AND intern(506) AND intern(507) AND intern(508) AND intern(509) AND intern(510) AND intern(511) AND intern(512)) OR ((NOT intern(505)) AND (NOT intern(506)) AND (NOT intern(507)) AND (NOT intern(508)) AND (NOT intern(509)) AND (NOT intern(510)) AND (NOT intern(511)) AND (NOT intern(512)));
--	intr_out(64) 	 <= 	 (intern(513) AND intern(514) AND intern(515) AND intern(516) AND intern(517) AND intern(518) AND intern(519) AND intern(520)) OR ((NOT intern(513)) AND (NOT intern(514)) AND (NOT intern(515)) AND (NOT intern(516)) AND (NOT intern(517)) AND (NOT intern(518)) AND (NOT intern(519)) AND (NOT intern(520)));
--	intr_out(65) 	 <= 	 (intern(521) AND intern(522) AND intern(523) AND intern(524) AND intern(525) AND intern(526) AND intern(527) AND intern(528)) OR ((NOT intern(521)) AND (NOT intern(522)) AND (NOT intern(523)) AND (NOT intern(524)) AND (NOT intern(525)) AND (NOT intern(526)) AND (NOT intern(527)) AND (NOT intern(528)));
--	intr_out(66) 	 <= 	 (intern(529) AND intern(530) AND intern(531) AND intern(532) AND intern(533) AND intern(534) AND intern(535) AND intern(536)) OR ((NOT intern(529)) AND (NOT intern(530)) AND (NOT intern(531)) AND (NOT intern(532)) AND (NOT intern(533)) AND (NOT intern(534)) AND (NOT intern(535)) AND (NOT intern(536)));
--	intr_out(67) 	 <= 	 (intern(537) AND intern(538) AND intern(539) AND intern(540) AND intern(541) AND intern(542) AND intern(543) AND intern(544)) OR ((NOT intern(537)) AND (NOT intern(538)) AND (NOT intern(539)) AND (NOT intern(540)) AND (NOT intern(541)) AND (NOT intern(542)) AND (NOT intern(543)) AND (NOT intern(544)));
--	intr_out(68) 	 <= 	 (intern(545) AND intern(546) AND intern(547) AND intern(548) AND intern(549) AND intern(550) AND intern(551) AND intern(552)) OR ((NOT intern(545)) AND (NOT intern(546)) AND (NOT intern(547)) AND (NOT intern(548)) AND (NOT intern(549)) AND (NOT intern(550)) AND (NOT intern(551)) AND (NOT intern(552)));
--	intr_out(69) 	 <= 	 (intern(553) AND intern(554) AND intern(555) AND intern(556) AND intern(557) AND intern(558) AND intern(559) AND intern(560)) OR ((NOT intern(553)) AND (NOT intern(554)) AND (NOT intern(555)) AND (NOT intern(556)) AND (NOT intern(557)) AND (NOT intern(558)) AND (NOT intern(559)) AND (NOT intern(560)));
--	intr_out(70) 	 <= 	 (intern(561) AND intern(562) AND intern(563) AND intern(564) AND intern(565) AND intern(566) AND intern(567) AND intern(568)) OR ((NOT intern(561)) AND (NOT intern(562)) AND (NOT intern(563)) AND (NOT intern(564)) AND (NOT intern(565)) AND (NOT intern(566)) AND (NOT intern(567)) AND (NOT intern(568)));
--	intr_out(71) 	 <= 	 (intern(569) AND intern(570) AND intern(571) AND intern(572) AND intern(573) AND intern(574) AND intern(575) AND intern(576)) OR ((NOT intern(569)) AND (NOT intern(570)) AND (NOT intern(571)) AND (NOT intern(572)) AND (NOT intern(573)) AND (NOT intern(574)) AND (NOT intern(575)) AND (NOT intern(576)));
--	intr_out(72) 	 <= 	 (intern(577) AND intern(578) AND intern(579) AND intern(580) AND intern(581) AND intern(582) AND intern(583) AND intern(584)) OR ((NOT intern(577)) AND (NOT intern(578)) AND (NOT intern(579)) AND (NOT intern(580)) AND (NOT intern(581)) AND (NOT intern(582)) AND (NOT intern(583)) AND (NOT intern(584)));
--	intr_out(73) 	 <= 	 (intern(585) AND intern(586) AND intern(587) AND intern(588) AND intern(589) AND intern(590) AND intern(591) AND intern(592)) OR ((NOT intern(585)) AND (NOT intern(586)) AND (NOT intern(587)) AND (NOT intern(588)) AND (NOT intern(589)) AND (NOT intern(590)) AND (NOT intern(591)) AND (NOT intern(592)));
--	intr_out(74) 	 <= 	 (intern(593) AND intern(594) AND intern(595) AND intern(596) AND intern(597) AND intern(598) AND intern(599) AND intern(600)) OR ((NOT intern(593)) AND (NOT intern(594)) AND (NOT intern(595)) AND (NOT intern(596)) AND (NOT intern(597)) AND (NOT intern(598)) AND (NOT intern(599)) AND (NOT intern(600)));
--	intr_out(75) 	 <= 	 (intern(601) AND intern(602) AND intern(603) AND intern(604) AND intern(605) AND intern(606) AND intern(607) AND intern(608)) OR ((NOT intern(601)) AND (NOT intern(602)) AND (NOT intern(603)) AND (NOT intern(604)) AND (NOT intern(605)) AND (NOT intern(606)) AND (NOT intern(607)) AND (NOT intern(608)));
--	intr_out(76) 	 <= 	 (intern(609) AND intern(610) AND intern(611) AND intern(612) AND intern(613) AND intern(614) AND intern(615) AND intern(616)) OR ((NOT intern(609)) AND (NOT intern(610)) AND (NOT intern(611)) AND (NOT intern(612)) AND (NOT intern(613)) AND (NOT intern(614)) AND (NOT intern(615)) AND (NOT intern(616)));
--	intr_out(77) 	 <= 	 (intern(617) AND intern(618) AND intern(619) AND intern(620) AND intern(621) AND intern(622) AND intern(623) AND intern(624)) OR ((NOT intern(617)) AND (NOT intern(618)) AND (NOT intern(619)) AND (NOT intern(620)) AND (NOT intern(621)) AND (NOT intern(622)) AND (NOT intern(623)) AND (NOT intern(624)));
--	intr_out(78) 	 <= 	 (intern(625) AND intern(626) AND intern(627) AND intern(628) AND intern(629) AND intern(630) AND intern(631) AND intern(632)) OR ((NOT intern(625)) AND (NOT intern(626)) AND (NOT intern(627)) AND (NOT intern(628)) AND (NOT intern(629)) AND (NOT intern(630)) AND (NOT intern(631)) AND (NOT intern(632)));
--	intr_out(79) 	 <= 	 (intern(633) AND intern(634) AND intern(635) AND intern(636) AND intern(637) AND intern(638) AND intern(639) AND intern(640)) OR ((NOT intern(633)) AND (NOT intern(634)) AND (NOT intern(635)) AND (NOT intern(636)) AND (NOT intern(637)) AND (NOT intern(638)) AND (NOT intern(639)) AND (NOT intern(640)));
--	intr_out(80) 	 <= 	 (intern(641) AND intern(642) AND intern(643) AND intern(644) AND intern(645) AND intern(646) AND intern(647) AND intern(648)) OR ((NOT intern(641)) AND (NOT intern(642)) AND (NOT intern(643)) AND (NOT intern(644)) AND (NOT intern(645)) AND (NOT intern(646)) AND (NOT intern(647)) AND (NOT intern(648)));
--	intr_out(81) 	 <= 	 (intern(649) AND intern(650) AND intern(651) AND intern(652) AND intern(653) AND intern(654) AND intern(655) AND intern(656)) OR ((NOT intern(649)) AND (NOT intern(650)) AND (NOT intern(651)) AND (NOT intern(652)) AND (NOT intern(653)) AND (NOT intern(654)) AND (NOT intern(655)) AND (NOT intern(656)));
--	intr_out(82) 	 <= 	 (intern(657) AND intern(658) AND intern(659) AND intern(660) AND intern(661) AND intern(662) AND intern(663) AND intern(664)) OR ((NOT intern(657)) AND (NOT intern(658)) AND (NOT intern(659)) AND (NOT intern(660)) AND (NOT intern(661)) AND (NOT intern(662)) AND (NOT intern(663)) AND (NOT intern(664)));
--	intr_out(83) 	 <= 	 (intern(665) AND intern(666) AND intern(667) AND intern(668) AND intern(669) AND intern(670) AND intern(671) AND intern(672)) OR ((NOT intern(665)) AND (NOT intern(666)) AND (NOT intern(667)) AND (NOT intern(668)) AND (NOT intern(669)) AND (NOT intern(670)) AND (NOT intern(671)) AND (NOT intern(672)));
--	intr_out(84) 	 <= 	 (intern(673) AND intern(674) AND intern(675) AND intern(676) AND intern(677) AND intern(678) AND intern(679) AND intern(680)) OR ((NOT intern(673)) AND (NOT intern(674)) AND (NOT intern(675)) AND (NOT intern(676)) AND (NOT intern(677)) AND (NOT intern(678)) AND (NOT intern(679)) AND (NOT intern(680)));
--	intr_out(85) 	 <= 	 (intern(681) AND intern(682) AND intern(683) AND intern(684) AND intern(685) AND intern(686) AND intern(687) AND intern(688)) OR ((NOT intern(681)) AND (NOT intern(682)) AND (NOT intern(683)) AND (NOT intern(684)) AND (NOT intern(685)) AND (NOT intern(686)) AND (NOT intern(687)) AND (NOT intern(688)));
--	intr_out(86) 	 <= 	 (intern(689) AND intern(690) AND intern(691) AND intern(692) AND intern(693) AND intern(694) AND intern(695) AND intern(696)) OR ((NOT intern(689)) AND (NOT intern(690)) AND (NOT intern(691)) AND (NOT intern(692)) AND (NOT intern(693)) AND (NOT intern(694)) AND (NOT intern(695)) AND (NOT intern(696)));
--	intr_out(87) 	 <= 	 (intern(697) AND intern(698) AND intern(699) AND intern(700) AND intern(701) AND intern(702) AND intern(703) AND intern(704)) OR ((NOT intern(697)) AND (NOT intern(698)) AND (NOT intern(699)) AND (NOT intern(700)) AND (NOT intern(701)) AND (NOT intern(702)) AND (NOT intern(703)) AND (NOT intern(704)));
--	intr_out(88) 	 <= 	 (intern(705) AND intern(706) AND intern(707) AND intern(708) AND intern(709) AND intern(710) AND intern(711) AND intern(712)) OR ((NOT intern(705)) AND (NOT intern(706)) AND (NOT intern(707)) AND (NOT intern(708)) AND (NOT intern(709)) AND (NOT intern(710)) AND (NOT intern(711)) AND (NOT intern(712)));
--	intr_out(89) 	 <= 	 (intern(713) AND intern(714) AND intern(715) AND intern(716) AND intern(717) AND intern(718) AND intern(719) AND intern(720)) OR ((NOT intern(713)) AND (NOT intern(714)) AND (NOT intern(715)) AND (NOT intern(716)) AND (NOT intern(717)) AND (NOT intern(718)) AND (NOT intern(719)) AND (NOT intern(720)));
--	intr_out(90) 	 <= 	 (intern(721) AND intern(722) AND intern(723) AND intern(724) AND intern(725) AND intern(726) AND intern(727) AND intern(728)) OR ((NOT intern(721)) AND (NOT intern(722)) AND (NOT intern(723)) AND (NOT intern(724)) AND (NOT intern(725)) AND (NOT intern(726)) AND (NOT intern(727)) AND (NOT intern(728)));
--	intr_out(91) 	 <= 	 (intern(729) AND intern(730) AND intern(731) AND intern(732) AND intern(733) AND intern(734) AND intern(735) AND intern(736)) OR ((NOT intern(729)) AND (NOT intern(730)) AND (NOT intern(731)) AND (NOT intern(732)) AND (NOT intern(733)) AND (NOT intern(734)) AND (NOT intern(735)) AND (NOT intern(736)));
--	intr_out(92) 	 <= 	 (intern(737) AND intern(738) AND intern(739) AND intern(740) AND intern(741) AND intern(742) AND intern(743) AND intern(744)) OR ((NOT intern(737)) AND (NOT intern(738)) AND (NOT intern(739)) AND (NOT intern(740)) AND (NOT intern(741)) AND (NOT intern(742)) AND (NOT intern(743)) AND (NOT intern(744)));
--	intr_out(93) 	 <= 	 (intern(745) AND intern(746) AND intern(747) AND intern(748) AND intern(749) AND intern(750) AND intern(751) AND intern(752)) OR ((NOT intern(745)) AND (NOT intern(746)) AND (NOT intern(747)) AND (NOT intern(748)) AND (NOT intern(749)) AND (NOT intern(750)) AND (NOT intern(751)) AND (NOT intern(752)));
--	intr_out(94) 	 <= 	 (intern(753) AND intern(754) AND intern(755) AND intern(756) AND intern(757) AND intern(758) AND intern(759) AND intern(760)) OR ((NOT intern(753)) AND (NOT intern(754)) AND (NOT intern(755)) AND (NOT intern(756)) AND (NOT intern(757)) AND (NOT intern(758)) AND (NOT intern(759)) AND (NOT intern(760)));
--	intr_out(95) 	 <= 	 (intern(761) AND intern(762) AND intern(763) AND intern(764) AND intern(765) AND intern(766) AND intern(767) AND intern(768)) OR ((NOT intern(761)) AND (NOT intern(762)) AND (NOT intern(763)) AND (NOT intern(764)) AND (NOT intern(765)) AND (NOT intern(766)) AND (NOT intern(767)) AND (NOT intern(768)));
--	intr_out(96) 	 <= 	 (intern(769) AND intern(770) AND intern(771) AND intern(772) AND intern(773) AND intern(774) AND intern(775) AND intern(776)) OR ((NOT intern(769)) AND (NOT intern(770)) AND (NOT intern(771)) AND (NOT intern(772)) AND (NOT intern(773)) AND (NOT intern(774)) AND (NOT intern(775)) AND (NOT intern(776)));
--	intr_out(97) 	 <= 	 (intern(777) AND intern(778) AND intern(779) AND intern(780) AND intern(781) AND intern(782) AND intern(783) AND intern(784)) OR ((NOT intern(777)) AND (NOT intern(778)) AND (NOT intern(779)) AND (NOT intern(780)) AND (NOT intern(781)) AND (NOT intern(782)) AND (NOT intern(783)) AND (NOT intern(784)));
--	intr_out(98) 	 <= 	 (intern(785) AND intern(786) AND intern(787) AND intern(788) AND intern(789) AND intern(790) AND intern(791) AND intern(792)) OR ((NOT intern(785)) AND (NOT intern(786)) AND (NOT intern(787)) AND (NOT intern(788)) AND (NOT intern(789)) AND (NOT intern(790)) AND (NOT intern(791)) AND (NOT intern(792)));
--	intr_out(99) 	 <= 	 (intern(793) AND intern(794) AND intern(795) AND intern(796) AND intern(797) AND intern(798) AND intern(799) AND intern(800)) OR ((NOT intern(793)) AND (NOT intern(794)) AND (NOT intern(795)) AND (NOT intern(796)) AND (NOT intern(797)) AND (NOT intern(798)) AND (NOT intern(799)) AND (NOT intern(800)));
--	intr_out(100) 	 <= 	 (intern(801) AND intern(802) AND intern(803) AND intern(804) AND intern(805) AND intern(806) AND intern(807) AND intern(808)) OR ((NOT intern(801)) AND (NOT intern(802)) AND (NOT intern(803)) AND (NOT intern(804)) AND (NOT intern(805)) AND (NOT intern(806)) AND (NOT intern(807)) AND (NOT intern(808)));
--	intr_out(101) 	 <= 	 (intern(809) AND intern(810) AND intern(811) AND intern(812) AND intern(813) AND intern(814) AND intern(815) AND intern(816)) OR ((NOT intern(809)) AND (NOT intern(810)) AND (NOT intern(811)) AND (NOT intern(812)) AND (NOT intern(813)) AND (NOT intern(814)) AND (NOT intern(815)) AND (NOT intern(816)));
--	intr_out(102) 	 <= 	 (intern(817) AND intern(818) AND intern(819) AND intern(820) AND intern(821) AND intern(822) AND intern(823) AND intern(824)) OR ((NOT intern(817)) AND (NOT intern(818)) AND (NOT intern(819)) AND (NOT intern(820)) AND (NOT intern(821)) AND (NOT intern(822)) AND (NOT intern(823)) AND (NOT intern(824)));
--	intr_out(103) 	 <= 	 (intern(825) AND intern(826) AND intern(827) AND intern(828) AND intern(829) AND intern(830) AND intern(831) AND intern(832)) OR ((NOT intern(825)) AND (NOT intern(826)) AND (NOT intern(827)) AND (NOT intern(828)) AND (NOT intern(829)) AND (NOT intern(830)) AND (NOT intern(831)) AND (NOT intern(832)));
--	intr_out(104) 	 <= 	 (intern(833) AND intern(834) AND intern(835) AND intern(836) AND intern(837) AND intern(838) AND intern(839) AND intern(840)) OR ((NOT intern(833)) AND (NOT intern(834)) AND (NOT intern(835)) AND (NOT intern(836)) AND (NOT intern(837)) AND (NOT intern(838)) AND (NOT intern(839)) AND (NOT intern(840)));
--	intr_out(105) 	 <= 	 (intern(841) AND intern(842) AND intern(843) AND intern(844) AND intern(845) AND intern(846) AND intern(847) AND intern(848)) OR ((NOT intern(841)) AND (NOT intern(842)) AND (NOT intern(843)) AND (NOT intern(844)) AND (NOT intern(845)) AND (NOT intern(846)) AND (NOT intern(847)) AND (NOT intern(848)));
--	intr_out(106) 	 <= 	 (intern(849) AND intern(850) AND intern(851) AND intern(852) AND intern(853) AND intern(854) AND intern(855) AND intern(856)) OR ((NOT intern(849)) AND (NOT intern(850)) AND (NOT intern(851)) AND (NOT intern(852)) AND (NOT intern(853)) AND (NOT intern(854)) AND (NOT intern(855)) AND (NOT intern(856)));
--	intr_out(107) 	 <= 	 (intern(857) AND intern(858) AND intern(859) AND intern(860) AND intern(861) AND intern(862) AND intern(863) AND intern(864)) OR ((NOT intern(857)) AND (NOT intern(858)) AND (NOT intern(859)) AND (NOT intern(860)) AND (NOT intern(861)) AND (NOT intern(862)) AND (NOT intern(863)) AND (NOT intern(864)));
--	intr_out(108) 	 <= 	 (intern(865) AND intern(866) AND intern(867) AND intern(868) AND intern(869) AND intern(870) AND intern(871) AND intern(872)) OR ((NOT intern(865)) AND (NOT intern(866)) AND (NOT intern(867)) AND (NOT intern(868)) AND (NOT intern(869)) AND (NOT intern(870)) AND (NOT intern(871)) AND (NOT intern(872)));
--	intr_out(109) 	 <= 	 (intern(873) AND intern(874) AND intern(875) AND intern(876) AND intern(877) AND intern(878) AND intern(879) AND intern(880)) OR ((NOT intern(873)) AND (NOT intern(874)) AND (NOT intern(875)) AND (NOT intern(876)) AND (NOT intern(877)) AND (NOT intern(878)) AND (NOT intern(879)) AND (NOT intern(880)));
--	intr_out(110) 	 <= 	 (intern(881) AND intern(882) AND intern(883) AND intern(884) AND intern(885) AND intern(886) AND intern(887) AND intern(888)) OR ((NOT intern(881)) AND (NOT intern(882)) AND (NOT intern(883)) AND (NOT intern(884)) AND (NOT intern(885)) AND (NOT intern(886)) AND (NOT intern(887)) AND (NOT intern(888)));
--	intr_out(111) 	 <= 	 (intern(889) AND intern(890) AND intern(891) AND intern(892) AND intern(893) AND intern(894) AND intern(895) AND intern(896)) OR ((NOT intern(889)) AND (NOT intern(890)) AND (NOT intern(891)) AND (NOT intern(892)) AND (NOT intern(893)) AND (NOT intern(894)) AND (NOT intern(895)) AND (NOT intern(896)));
--	intr_out(112) 	 <= 	 (intern(897) AND intern(898) AND intern(899) AND intern(900) AND intern(901) AND intern(902) AND intern(903) AND intern(904)) OR ((NOT intern(897)) AND (NOT intern(898)) AND (NOT intern(899)) AND (NOT intern(900)) AND (NOT intern(901)) AND (NOT intern(902)) AND (NOT intern(903)) AND (NOT intern(904)));
--	intr_out(113) 	 <= 	 (intern(905) AND intern(906) AND intern(907) AND intern(908) AND intern(909) AND intern(910) AND intern(911) AND intern(912)) OR ((NOT intern(905)) AND (NOT intern(906)) AND (NOT intern(907)) AND (NOT intern(908)) AND (NOT intern(909)) AND (NOT intern(910)) AND (NOT intern(911)) AND (NOT intern(912)));
--	intr_out(114) 	 <= 	 (intern(913) AND intern(914) AND intern(915) AND intern(916) AND intern(917) AND intern(918) AND intern(919) AND intern(920)) OR ((NOT intern(913)) AND (NOT intern(914)) AND (NOT intern(915)) AND (NOT intern(916)) AND (NOT intern(917)) AND (NOT intern(918)) AND (NOT intern(919)) AND (NOT intern(920)));
--	intr_out(115) 	 <= 	 (intern(921) AND intern(922) AND intern(923) AND intern(924) AND intern(925) AND intern(926) AND intern(927) AND intern(928)) OR ((NOT intern(921)) AND (NOT intern(922)) AND (NOT intern(923)) AND (NOT intern(924)) AND (NOT intern(925)) AND (NOT intern(926)) AND (NOT intern(927)) AND (NOT intern(928)));
--	intr_out(116) 	 <= 	 (intern(929) AND intern(930) AND intern(931) AND intern(932) AND intern(933) AND intern(934) AND intern(935) AND intern(936)) OR ((NOT intern(929)) AND (NOT intern(930)) AND (NOT intern(931)) AND (NOT intern(932)) AND (NOT intern(933)) AND (NOT intern(934)) AND (NOT intern(935)) AND (NOT intern(936)));
--	intr_out(117) 	 <= 	 (intern(937) AND intern(938) AND intern(939) AND intern(940) AND intern(941) AND intern(942) AND intern(943) AND intern(944)) OR ((NOT intern(937)) AND (NOT intern(938)) AND (NOT intern(939)) AND (NOT intern(940)) AND (NOT intern(941)) AND (NOT intern(942)) AND (NOT intern(943)) AND (NOT intern(944)));
--	intr_out(118) 	 <= 	 (intern(945) AND intern(946) AND intern(947) AND intern(948) AND intern(949) AND intern(950) AND intern(951) AND intern(952)) OR ((NOT intern(945)) AND (NOT intern(946)) AND (NOT intern(947)) AND (NOT intern(948)) AND (NOT intern(949)) AND (NOT intern(950)) AND (NOT intern(951)) AND (NOT intern(952)));
--	intr_out(119) 	 <= 	 (intern(953) AND intern(954) AND intern(955) AND intern(956) AND intern(957) AND intern(958) AND intern(959) AND intern(960)) OR ((NOT intern(953)) AND (NOT intern(954)) AND (NOT intern(955)) AND (NOT intern(956)) AND (NOT intern(957)) AND (NOT intern(958)) AND (NOT intern(959)) AND (NOT intern(960)));
--	intr_out(120) 	 <= 	 (intern(961) AND intern(962) AND intern(963) AND intern(964) AND intern(965) AND intern(966) AND intern(967) AND intern(968)) OR ((NOT intern(961)) AND (NOT intern(962)) AND (NOT intern(963)) AND (NOT intern(964)) AND (NOT intern(965)) AND (NOT intern(966)) AND (NOT intern(967)) AND (NOT intern(968)));
--	intr_out(121) 	 <= 	 (intern(969) AND intern(970) AND intern(971) AND intern(972) AND intern(973) AND intern(974) AND intern(975) AND intern(976)) OR ((NOT intern(969)) AND (NOT intern(970)) AND (NOT intern(971)) AND (NOT intern(972)) AND (NOT intern(973)) AND (NOT intern(974)) AND (NOT intern(975)) AND (NOT intern(976)));
--	intr_out(122) 	 <= 	 (intern(977) AND intern(978) AND intern(979) AND intern(980) AND intern(981) AND intern(982) AND intern(983) AND intern(984)) OR ((NOT intern(977)) AND (NOT intern(978)) AND (NOT intern(979)) AND (NOT intern(980)) AND (NOT intern(981)) AND (NOT intern(982)) AND (NOT intern(983)) AND (NOT intern(984)));
--	intr_out(123) 	 <= 	 (intern(985) AND intern(986) AND intern(987) AND intern(988) AND intern(989) AND intern(990) AND intern(991) AND intern(992)) OR ((NOT intern(985)) AND (NOT intern(986)) AND (NOT intern(987)) AND (NOT intern(988)) AND (NOT intern(989)) AND (NOT intern(990)) AND (NOT intern(991)) AND (NOT intern(992)));
--	intr_out(124) 	 <= 	 (intern(993) AND intern(994) AND intern(995) AND intern(996) AND intern(997) AND intern(998) AND intern(999) AND intern(1000)) OR ((NOT intern(993)) AND (NOT intern(994)) AND (NOT intern(995)) AND (NOT intern(996)) AND (NOT intern(997)) AND (NOT intern(998)) AND (NOT intern(999)) AND (NOT intern(1000)));
--	intr_out(125) 	 <= 	 (intern(1001) AND intern(1002) AND intern(1003) AND intern(1004) AND intern(1005) AND intern(1006) AND intern(1007) AND intern(1008)) OR ((NOT intern(1001)) AND (NOT intern(1002)) AND (NOT intern(1003)) AND (NOT intern(1004)) AND (NOT intern(1005)) AND (NOT intern(1006)) AND (NOT intern(1007)) AND (NOT intern(1008)));
--	intr_out(126) 	 <= 	 (intern(1009) AND intern(1010) AND intern(1011) AND intern(1012) AND intern(1013) AND intern(1014) AND intern(1015) AND intern(1016)) OR ((NOT intern(1009)) AND (NOT intern(1010)) AND (NOT intern(1011)) AND (NOT intern(1012)) AND (NOT intern(1013)) AND (NOT intern(1014)) AND (NOT intern(1015)) AND (NOT intern(1016)));
--	intr_out(127) 	 <= 	 (intern(1017) AND intern(1018) AND intern(1019) AND intern(1020) AND intern(1021) AND intern(1022) AND intern(1023)) OR ((NOT intern(1017)) AND (NOT intern(1018)) AND (NOT intern(1019)) AND (NOT intern(1020)) AND (NOT intern(1021)) AND (NOT intern(1022)) AND (NOT intern(1023)));

	reset <= rst;
	
end structural ;

